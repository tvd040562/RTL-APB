VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO apb_memory
  CLASS BLOCK ;
  FOREIGN apb_memory ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN paddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END paddr[0]
  PIN paddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END paddr[1]
  PIN paddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END paddr[2]
  PIN paddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END paddr[3]
  PIN pclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END pclk
  PIN prdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 54.440 150.000 55.040 ;
    END
  END prdata[0]
  PIN prdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 44.240 150.000 44.840 ;
    END
  END prdata[1]
  PIN prdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.240 150.000 78.840 ;
    END
  END prdata[2]
  PIN prdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.040 150.000 68.640 ;
    END
  END prdata[3]
  PIN prdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 51.040 150.000 51.640 ;
    END
  END prdata[4]
  PIN prdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 64.640 150.000 65.240 ;
    END
  END prdata[5]
  PIN prdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.840 150.000 75.440 ;
    END
  END prdata[6]
  PIN prdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 71.440 150.000 72.040 ;
    END
  END prdata[7]
  PIN pwdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END pwdata[0]
  PIN pwdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END pwdata[1]
  PIN pwdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END pwdata[2]
  PIN pwdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END pwdata[3]
  PIN pwdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END pwdata[4]
  PIN pwdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 146.000 84.090 150.000 ;
    END
  END pwdata[5]
  PIN pwdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END pwdata[6]
  PIN pwdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END pwdata[7]
  PIN ren
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 61.240 150.000 61.840 ;
    END
  END ren
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 47.640 150.000 48.240 ;
    END
  END rst_n
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 138.960 ;
    END
  END vssd1
  PIN wen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 57.840 150.000 58.440 ;
    END
  END wen
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 4.670 10.640 144.830 138.960 ;
      LAYER met2 ;
        RECT 4.690 145.720 83.530 146.610 ;
        RECT 84.370 145.720 144.810 146.610 ;
        RECT 4.690 4.280 144.810 145.720 ;
        RECT 4.690 4.000 41.670 4.280 ;
        RECT 42.510 4.000 54.550 4.280 ;
        RECT 55.390 4.000 144.810 4.280 ;
      LAYER met3 ;
        RECT 3.990 137.040 146.000 138.885 ;
        RECT 4.400 135.640 146.000 137.040 ;
        RECT 3.990 133.640 146.000 135.640 ;
        RECT 4.400 132.240 146.000 133.640 ;
        RECT 3.990 123.440 146.000 132.240 ;
        RECT 4.400 122.040 146.000 123.440 ;
        RECT 3.990 120.040 146.000 122.040 ;
        RECT 4.400 118.640 146.000 120.040 ;
        RECT 3.990 116.640 146.000 118.640 ;
        RECT 4.400 115.240 146.000 116.640 ;
        RECT 3.990 99.640 146.000 115.240 ;
        RECT 4.400 98.240 146.000 99.640 ;
        RECT 3.990 86.040 146.000 98.240 ;
        RECT 4.400 84.640 146.000 86.040 ;
        RECT 3.990 82.640 146.000 84.640 ;
        RECT 4.400 81.240 146.000 82.640 ;
        RECT 3.990 79.240 146.000 81.240 ;
        RECT 4.400 77.840 145.600 79.240 ;
        RECT 3.990 75.840 146.000 77.840 ;
        RECT 4.400 74.440 145.600 75.840 ;
        RECT 3.990 72.440 146.000 74.440 ;
        RECT 4.400 71.040 145.600 72.440 ;
        RECT 3.990 69.040 146.000 71.040 ;
        RECT 4.400 67.640 145.600 69.040 ;
        RECT 3.990 65.640 146.000 67.640 ;
        RECT 3.990 64.240 145.600 65.640 ;
        RECT 3.990 62.240 146.000 64.240 ;
        RECT 3.990 60.840 145.600 62.240 ;
        RECT 3.990 58.840 146.000 60.840 ;
        RECT 3.990 57.440 145.600 58.840 ;
        RECT 3.990 55.440 146.000 57.440 ;
        RECT 3.990 54.040 145.600 55.440 ;
        RECT 3.990 52.040 146.000 54.040 ;
        RECT 3.990 50.640 145.600 52.040 ;
        RECT 3.990 48.640 146.000 50.640 ;
        RECT 3.990 47.240 145.600 48.640 ;
        RECT 3.990 45.240 146.000 47.240 ;
        RECT 3.990 43.840 145.600 45.240 ;
        RECT 3.990 10.715 146.000 43.840 ;
      LAYER met4 ;
        RECT 110.695 47.775 123.905 103.865 ;
  END
END apb_memory
END LIBRARY

